library IEEE;
use IEEE.STD_LOGIC_1164.all;

package CONSTANTS is 
	constant NumBit 			: integer := 14;
	constant Nt 				: integer := 8;
	constant shift				: integer := 7;
    constant MAX_DEC    		: integer := 8192;
	constant unfolding_stages 	: integer := 3;
end CONSTANTS;
